module fetch_cycle(clk,rst,);