module Controller(instr,RegWE);

input [31:0]instr;
output RegWE;

