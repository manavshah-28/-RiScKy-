/*/////////////////////////////////////////////
 File: Regfile.v
 Author: Manav Shah
 ----------------------------------------------

    ██████╗ ██╗███████╗ ██████╗██╗  ██╗██╗   ██╗
    ██╔══██╗██║██╔════╝██╔════╝██║ ██╔╝╚██╗ ██╔╝
    ██████╔╝██║███████╗██║     █████╔╝  ╚████╔╝ 
    ██╔══██╗██║╚════██║██║     ██╔═██╗   ╚██╔╝  
    ██║  ██║██║███████║╚██████╗██║  ██╗   ██║   
    ╚═╝  ╚═╝╚═╝╚══════╝ ╚═════╝╚═╝  ╚═╝   ╚═╝   
 ----------------------------------------------
                                    
 Copyright (c) 2024 MANAV SHAH
*//////////////////////////////////////////////

module Regfile(clk,rst,WE,AddD,DataD,AddA,DataA,AddB,DataB);
input clk,rst,WE;
input [4:0] AddA,AddB,AddD;
input [31:0] DataD;
/*
rst: is reset signal(active low).
WE: is Write Enable signal.
AddA,AddB : registers are read at these addresses
and read values are given out at DataA and DataB respectively.
AddD : is the address for the register which is to be written with DataD.
*/
output [31:0] DataA,DataB;

logic [31:0] xreg [31:0]; //x0 to x31 : RV32 registers
logic [4:0]index = 1;

initial begin
foreach (xreg[i]) begin
    xreg[i] = 'd0;
end
end
// initial begin
//     $readmemh("reg_load.hex",xreg,0,31); // custom program to load registers from gui
// end

always @(posedge clk)begin
   if(WE &(AddD != 5'h00))
       xreg[AddD] <= DataD;  
end

assign DataA = (rst == 1'b0) ? 32'h00000000 : xreg[AddA];
assign DataB = (rst == 1'b0) ? 32'h00000000 : xreg[AddB];

endmodule

