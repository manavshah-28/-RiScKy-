module branch_comp(A,B,BrUn,BrEq,BrLt);

input [31:0]A,B;
input BrUn;

output BrEq,BrLt;

endmodule